.subckt comparator N001 N002 0 N006 N005 Vout
M1 N003 N003 N001 N001 pfet l=200n w=2u m=1
M2 N004 N003 N001 N001 pfet l=200n w=2u m=1
M3 N003 N005 N008 0 nfet l=200n w=2u m=1
M4 N004 N006 N008 0 nfet l=200n w=2u m=1
M5 N009 N004 N001 N001 pfet l=200n w=6u m=1
M6 N009 N007 0 0 nfet l=200n w=2u m=1
M7 N008 N007 0 0 nfet l=200n w=2u m=1
M8 N010 N009 N002 N002 pfet l=200n w=2u
M9 Vout N010 N002 N002 pfet l=200n w=2u
M10 N010 N009 0 0 nfet l=200n w=1u
M11 Vout N010 0 0 nfet l=200n w=1u
*C1 Vout 0 1f
*C2 N009 0 1f
*M12 N007 clk N001 N001 pfet l=0.2u w=3u
*I1 N001 N007 2u
R N001 N007 10k
M13 N007 N007 0 0 nfet l=0.2u w=2u
.ends comparator


X1 1 1d 0 v_p v_n out_comp comparator

V_a 1 0 3.3v
V_d 1d 0 1.8V


Vp v_p 0 pulse(2.06 0 1n 1n 1n 1u 2u)
Vn v_n 0 pulse(0 2.06 1n 1n 1n 1u 2u)
